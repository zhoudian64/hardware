module ascii(
    input   [31:0]  program_counter,
    output  [31:0]  instruction,
);
wire   [31:0] rom [0:63];
assign rom[6'h00] = 32'b11000000000000000000100100110111; //
assign rom[6'h01] = 32'b10100000000000000000100110110111; //
assign rom[6'h02] = 32'b00000000000000000000001010010011; //
assign rom[6'h03] = 32'b00000000000000000000001100010011; //
assign rom[6'h04] = 32'b00000101000000000000011010010011; //
assign rom[6'h05] = 32'b11111111111111110000011100110111; //
assign rom[6'h06] = 32'b00000000111010011010000000100011; //
assign rom[6'h07] = 32'b00000000000010011010010100000011; //
assign rom[6'h08] = 32'b00010000000001010111010110010011; //
assign rom[6'h09] = 32'b11111110000001011000110011100011; //
assign rom[6'h0a] = 32'b00001111111101010111010110010011; //
assign rom[6'h0b] = 32'b00000000010001011101010100010011; //
assign rom[6'h0c] = 32'b00000010000000000000000011101111; //
assign rom[6'h0d] = 32'b00000011010000000000000011101111; //
assign rom[6'h0e] = 32'b00000000111101011111010100010011; //
assign rom[6'h0f] = 32'b00000001010000000000000011101111; //
assign rom[6'h10] = 32'b00000010100000000000000011101111; //
assign rom[6'h11] = 32'b00000010000000000000010100010011; //
assign rom[6'h12] = 32'b00000010000000000000000011101111; //
assign rom[6'h13] = 32'b11111101000111111111000001101111; //
assign rom[6'h14] = 32'b11111111011101010000001110010011; //
assign rom[6'h15] = 32'b00000000011100000100011001100011; //
assign rom[6'h16] = 32'b00000011000001010000010100010011; //
assign rom[6'h17] = 32'b00000000000000001000000001100111; //
assign rom[6'h18] = 32'b00000011011101010000010100010011; //
assign rom[6'h19] = 32'b00000000000000001000000001100111; //
assign rom[6'h1a] = 32'b00000000101010010010000000100011; //
assign rom[6'h1b] = 32'b00000000010010010000100100010011; //
assign rom[6'h1c] = 32'b00000000000100110000001100010011; //
assign rom[6'h1d] = 32'b00000000110100110001011001100011; //
assign rom[6'h1e] = 32'b00000000000100101000001010010011; //
assign rom[6'h1f] = 32'b00000000000000000000001100010011; //
assign rom[6'h20] = 32'b00000000100000101001111000010011; //
assign rom[6'h21] = 32'b00000000011011100110111000110011; //
assign rom[6'h22] = 32'b11111111111111110000011100110111; //
assign rom[6'h23] = 32'b00000001110001110110011100110011; //
assign rom[6'h24] = 32'b00000000111010011010000000100011; //
assign rom[6'h25] = 32'b00000000000000001000000001100111; //
assign rom[6'h26] = 32'b00000000000000000000000000000000; //
assign rom[6'h27] = 32'b00000000000000000000000000000000; //
assign rom[6'h28] = 32'b00000000000000000000000000000000; //
assign rom[6'h29] = 32'b00000000000000000000000000000000; //
assign rom[6'h2a] = 32'b00000000000000000000000000000000; //
assign rom[6'h2b] = 32'b00000000000000000000000000000000; //
assign rom[6'h2c] = 32'b00000000000000000000000000000000; //
assign rom[6'h2d] = 32'b00000000000000000000000000000000; //
assign rom[6'h2e] = 32'b00000000000000000000000000000000; //
assign rom[6'h2f] = 32'b00000000000000000000000000000000; //
assign rom[6'h30] = 32'b00000000000000000000000000000000; //
assign rom[6'h31] = 32'b00000000000000000000000000000000; //
assign rom[6'h32] = 32'b00000000000000000000000000000000; //
assign rom[6'h33] = 32'b00000000000000000000000000000000; //
assign rom[6'h34] = 32'b00000000000000000000000000000000; //
assign rom[6'h35] = 32'b00000000000000000000000000000000; //
assign rom[6'h36] = 32'b00000000000000000000000000000000; //
assign rom[6'h37] = 32'b00000000000000000000000000000000; //
assign rom[6'h38] = 32'b00000000000000000000000000000000; //
assign rom[6'h39] = 32'b00000000000000000000000000000000; //
assign rom[6'h3a] = 32'b00000000000000000000000000000000; //
assign rom[6'h3b] = 32'b00000000000000000000000000000000; //
assign rom[6'h3c] = 32'b00000000000000000000000000000000; //
assign rom[6'h3d] = 32'b00000000000000000000000000000000; //
assign rom[6'h3e] = 32'b00000000000000000000000000000000; //
assign rom[6'h3f] = 32'b00000000000000000000000000000000; //
assign instruction = rom[program_counter[7:2]];

endmodule // ascii.v